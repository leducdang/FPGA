// I2C.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module I2C (
		input  wire  clk_clk,       //   clk.clk
		input  wire  i2c_sda_in,    //   i2c.sda_in
		input  wire  i2c_scl_in,    //      .scl_in
		output wire  i2c_sda_oe,    //      .sda_oe
		output wire  i2c_scl_oe,    //      .scl_oe
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire  [31:0] cpu_data_master_readdata;                              // mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_waitrequest;                           // mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire         cpu_data_master_debugaccess;                           // CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	wire  [19:0] cpu_data_master_address;                               // CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                            // CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	wire         cpu_data_master_read;                                  // CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	wire         cpu_data_master_write;                                 // CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	wire  [31:0] cpu_data_master_writedata;                             // CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                       // mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_waitrequest;                    // mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [19:0] cpu_instruction_master_address;                        // CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                           // CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	wire         mm_interconnect_0_debug_avalon_jtag_slave_chipselect;  // mm_interconnect_0:DEBUG_avalon_jtag_slave_chipselect -> DEBUG:av_chipselect
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_readdata;    // DEBUG:av_readdata -> mm_interconnect_0:DEBUG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_debug_avalon_jtag_slave_waitrequest; // DEBUG:av_waitrequest -> mm_interconnect_0:DEBUG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_debug_avalon_jtag_slave_address;     // mm_interconnect_0:DEBUG_avalon_jtag_slave_address -> DEBUG:av_address
	wire         mm_interconnect_0_debug_avalon_jtag_slave_read;        // mm_interconnect_0:DEBUG_avalon_jtag_slave_read -> DEBUG:av_read_n
	wire         mm_interconnect_0_debug_avalon_jtag_slave_write;       // mm_interconnect_0:DEBUG_avalon_jtag_slave_write -> DEBUG:av_write_n
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_writedata;   // mm_interconnect_0:DEBUG_avalon_jtag_slave_writedata -> DEBUG:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata; // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;  // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_i2c_csr_readdata;                    // I2C:readdata -> mm_interconnect_0:I2C_csr_readdata
	wire   [3:0] mm_interconnect_0_i2c_csr_address;                     // mm_interconnect_0:I2C_csr_address -> I2C:addr
	wire         mm_interconnect_0_i2c_csr_read;                        // mm_interconnect_0:I2C_csr_read -> I2C:read
	wire         mm_interconnect_0_i2c_csr_write;                       // mm_interconnect_0:I2C_csr_write -> I2C:write
	wire  [31:0] mm_interconnect_0_i2c_csr_writedata;                   // mm_interconnect_0:I2C_csr_writedata -> I2C:writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;        // CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;     // CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;     // mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;         // mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;            // mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;      // mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;           // mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;       // mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                   // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                     // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [15:0] mm_interconnect_0_ram_s1_address;                      // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                   // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                        // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                    // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                        // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         mm_interconnect_0_timer_0_s1_chipselect;               // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                 // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                  // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                    // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         irq_mapper_receiver0_irq;                              // I2C:intr -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                              // DEBUG:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                              // timer_0:irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu_irq_irq;                                           // irq_mapper:sender_irq -> CPU:irq
	wire         rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [CPU:reset_n, DEBUG:rst_n, I2C:rst_n, RAM:reset, irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, sysid_qsys_0:reset_n, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                    // rst_controller:reset_req -> [CPU:reset_req, RAM:reset_req, rst_translator:reset_req_in]

	I2C_CPU cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	I2C_DEBUG debug (
		.clk            (clk_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_debug_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_debug_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_debug_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                               //               irq.irq
	);

	altera_avalon_i2c #(
		.USE_AV_ST       (0),
		.FIFO_DEPTH      (4),
		.FIFO_DEPTH_LOG2 (2)
	) i2c (
		.clk       (clk_clk),                             //            clock.clk
		.rst_n     (~rst_controller_reset_out_reset),     //       reset_sink.reset_n
		.intr      (irq_mapper_receiver0_irq),            // interrupt_sender.irq
		.addr      (mm_interconnect_0_i2c_csr_address),   //              csr.address
		.read      (mm_interconnect_0_i2c_csr_read),      //                 .read
		.write     (mm_interconnect_0_i2c_csr_write),     //                 .write
		.writedata (mm_interconnect_0_i2c_csr_writedata), //                 .writedata
		.readdata  (mm_interconnect_0_i2c_csr_readdata),  //                 .readdata
		.sda_in    (i2c_sda_in),                          //       i2c_serial.sda_in
		.scl_in    (i2c_scl_in),                          //                 .scl_in
		.sda_oe    (i2c_sda_oe),                          //                 .sda_oe
		.scl_oe    (i2c_scl_oe),                          //                 .scl_oe
		.src_data  (),                                    //      (terminated)
		.src_valid (),                                    //      (terminated)
		.src_ready (1'b0),                                //      (terminated)
		.snk_data  (16'b0000000000000000),                //      (terminated)
		.snk_valid (1'b0),                                //      (terminated)
		.snk_ready ()                                     //      (terminated)
	);

	I2C_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	I2C_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	I2C_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                 //   irq.irq
	);

	I2C_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                         (clk_clk),                                               //                       clk_0_clk.clk
		.CPU_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                        // CPU_reset_reset_bridge_in_reset.reset
		.CPU_data_master_address               (cpu_data_master_address),                               //                 CPU_data_master.address
		.CPU_data_master_waitrequest           (cpu_data_master_waitrequest),                           //                                .waitrequest
		.CPU_data_master_byteenable            (cpu_data_master_byteenable),                            //                                .byteenable
		.CPU_data_master_read                  (cpu_data_master_read),                                  //                                .read
		.CPU_data_master_readdata              (cpu_data_master_readdata),                              //                                .readdata
		.CPU_data_master_write                 (cpu_data_master_write),                                 //                                .write
		.CPU_data_master_writedata             (cpu_data_master_writedata),                             //                                .writedata
		.CPU_data_master_debugaccess           (cpu_data_master_debugaccess),                           //                                .debugaccess
		.CPU_instruction_master_address        (cpu_instruction_master_address),                        //          CPU_instruction_master.address
		.CPU_instruction_master_waitrequest    (cpu_instruction_master_waitrequest),                    //                                .waitrequest
		.CPU_instruction_master_read           (cpu_instruction_master_read),                           //                                .read
		.CPU_instruction_master_readdata       (cpu_instruction_master_readdata),                       //                                .readdata
		.CPU_debug_mem_slave_address           (mm_interconnect_0_cpu_debug_mem_slave_address),         //             CPU_debug_mem_slave.address
		.CPU_debug_mem_slave_write             (mm_interconnect_0_cpu_debug_mem_slave_write),           //                                .write
		.CPU_debug_mem_slave_read              (mm_interconnect_0_cpu_debug_mem_slave_read),            //                                .read
		.CPU_debug_mem_slave_readdata          (mm_interconnect_0_cpu_debug_mem_slave_readdata),        //                                .readdata
		.CPU_debug_mem_slave_writedata         (mm_interconnect_0_cpu_debug_mem_slave_writedata),       //                                .writedata
		.CPU_debug_mem_slave_byteenable        (mm_interconnect_0_cpu_debug_mem_slave_byteenable),      //                                .byteenable
		.CPU_debug_mem_slave_waitrequest       (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),     //                                .waitrequest
		.CPU_debug_mem_slave_debugaccess       (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),     //                                .debugaccess
		.DEBUG_avalon_jtag_slave_address       (mm_interconnect_0_debug_avalon_jtag_slave_address),     //         DEBUG_avalon_jtag_slave.address
		.DEBUG_avalon_jtag_slave_write         (mm_interconnect_0_debug_avalon_jtag_slave_write),       //                                .write
		.DEBUG_avalon_jtag_slave_read          (mm_interconnect_0_debug_avalon_jtag_slave_read),        //                                .read
		.DEBUG_avalon_jtag_slave_readdata      (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                                .readdata
		.DEBUG_avalon_jtag_slave_writedata     (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                                .writedata
		.DEBUG_avalon_jtag_slave_waitrequest   (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                                .waitrequest
		.DEBUG_avalon_jtag_slave_chipselect    (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  //                                .chipselect
		.I2C_csr_address                       (mm_interconnect_0_i2c_csr_address),                     //                         I2C_csr.address
		.I2C_csr_write                         (mm_interconnect_0_i2c_csr_write),                       //                                .write
		.I2C_csr_read                          (mm_interconnect_0_i2c_csr_read),                        //                                .read
		.I2C_csr_readdata                      (mm_interconnect_0_i2c_csr_readdata),                    //                                .readdata
		.I2C_csr_writedata                     (mm_interconnect_0_i2c_csr_writedata),                   //                                .writedata
		.RAM_s1_address                        (mm_interconnect_0_ram_s1_address),                      //                          RAM_s1.address
		.RAM_s1_write                          (mm_interconnect_0_ram_s1_write),                        //                                .write
		.RAM_s1_readdata                       (mm_interconnect_0_ram_s1_readdata),                     //                                .readdata
		.RAM_s1_writedata                      (mm_interconnect_0_ram_s1_writedata),                    //                                .writedata
		.RAM_s1_byteenable                     (mm_interconnect_0_ram_s1_byteenable),                   //                                .byteenable
		.RAM_s1_chipselect                     (mm_interconnect_0_ram_s1_chipselect),                   //                                .chipselect
		.RAM_s1_clken                          (mm_interconnect_0_ram_s1_clken),                        //                                .clken
		.sysid_qsys_0_control_slave_address    (mm_interconnect_0_sysid_qsys_0_control_slave_address),  //      sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata   (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), //                                .readdata
		.timer_0_s1_address                    (mm_interconnect_0_timer_0_s1_address),                  //                      timer_0_s1.address
		.timer_0_s1_write                      (mm_interconnect_0_timer_0_s1_write),                    //                                .write
		.timer_0_s1_readdata                   (mm_interconnect_0_timer_0_s1_readdata),                 //                                .readdata
		.timer_0_s1_writedata                  (mm_interconnect_0_timer_0_s1_writedata),                //                                .writedata
		.timer_0_s1_chipselect                 (mm_interconnect_0_timer_0_s1_chipselect)                //                                .chipselect
	);

	I2C_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
