
module step (
	clk_clk,
	reset_reset_n,
	out1_export,
	out2_export,
	out3_export,
	out4_export);	

	input		clk_clk;
	input		reset_reset_n;
	output		out1_export;
	output		out2_export;
	output		out3_export;
	output		out4_export;
endmodule
