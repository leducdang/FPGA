
module bai1 (
	clk_clk,
	led_export,
	reset_reset_n,
	bt1_export);	

	input		clk_clk;
	output	[7:0]	led_export;
	input		reset_reset_n;
	input		bt1_export;
endmodule
