
module ledMatrix (
	clk_clk,
	reset_reset_n,
	r1_export,
	r2_export,
	r3_export,
	r4_export,
	c1_export,
	c2_export,
	c3_export,
	c4_export);	

	input		clk_clk;
	input		reset_reset_n;
	output		r1_export;
	output		r2_export;
	output		r3_export;
	output		r4_export;
	input		c1_export;
	input		c2_export;
	input		c3_export;
	input		c4_export;
endmodule
