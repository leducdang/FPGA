module top(
				clock_50mhz,
				pin_reset,
				);
				

				
				
				
endmodule