// ed_sim.v

// Generated using ACDS version 22.1 915

`timescale 1 ps / 1 ps
module ed_sim (
		output wire [15:0] tg_pnf_pnf_per_bit,         // tg_pnf.pnf_per_bit
		output wire [15:0] tg_pnf_pnf_per_bit_persist  //       .pnf_per_bit_persist
	);

	ed_sim_ed_sim ed_sim (
		.tg_pnf_pnf_per_bit         (tg_pnf_pnf_per_bit),         // tg_pnf.pnf_per_bit
		.tg_pnf_pnf_per_bit_persist (tg_pnf_pnf_per_bit_persist)  //       .pnf_per_bit_persist
	);

endmodule
