
module bluetooth (
	clk_clk,
	reset_reset_n,
	rs232_RXD,
	rs232_TXD);	

	input		clk_clk;
	input		reset_reset_n;
	input		rs232_RXD;
	output		rs232_TXD;
endmodule
