// ledMatrix.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module ledMatrix (
		input  wire  c1_export,     //    c1.export
		input  wire  c2_export,     //    c2.export
		input  wire  c3_export,     //    c3.export
		input  wire  c4_export,     //    c4.export
		input  wire  clk_clk,       //   clk.clk
		output wire  r1_export,     //    r1.export
		output wire  r2_export,     //    r2.export
		output wire  r3_export,     //    r3.export
		output wire  r4_export,     //    r4.export
		input  wire  reset_reset_n  // reset.reset_n
	);

	wire  [31:0] cpu_data_master_readdata;                              // mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_waitrequest;                           // mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire         cpu_data_master_debugaccess;                           // CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	wire  [19:0] cpu_data_master_address;                               // CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                            // CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	wire         cpu_data_master_read;                                  // CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	wire         cpu_data_master_write;                                 // CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	wire  [31:0] cpu_data_master_writedata;                             // CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                       // mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_waitrequest;                    // mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [19:0] cpu_instruction_master_address;                        // CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                           // CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	wire         mm_interconnect_0_debug_avalon_jtag_slave_chipselect;  // mm_interconnect_0:DEBUG_avalon_jtag_slave_chipselect -> DEBUG:av_chipselect
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_readdata;    // DEBUG:av_readdata -> mm_interconnect_0:DEBUG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_debug_avalon_jtag_slave_waitrequest; // DEBUG:av_waitrequest -> mm_interconnect_0:DEBUG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_debug_avalon_jtag_slave_address;     // mm_interconnect_0:DEBUG_avalon_jtag_slave_address -> DEBUG:av_address
	wire         mm_interconnect_0_debug_avalon_jtag_slave_read;        // mm_interconnect_0:DEBUG_avalon_jtag_slave_read -> DEBUG:av_read_n
	wire         mm_interconnect_0_debug_avalon_jtag_slave_write;       // mm_interconnect_0:DEBUG_avalon_jtag_slave_write -> DEBUG:av_write_n
	wire  [31:0] mm_interconnect_0_debug_avalon_jtag_slave_writedata;   // mm_interconnect_0:DEBUG_avalon_jtag_slave_writedata -> DEBUG:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;        // CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;     // CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;     // mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;         // mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;            // mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;      // mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;           // mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;       // mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_c4_s1_readdata;                      // C4:readdata -> mm_interconnect_0:C4_s1_readdata
	wire   [1:0] mm_interconnect_0_c4_s1_address;                       // mm_interconnect_0:C4_s1_address -> C4:address
	wire  [31:0] mm_interconnect_0_c3_s1_readdata;                      // C3:readdata -> mm_interconnect_0:C3_s1_readdata
	wire   [1:0] mm_interconnect_0_c3_s1_address;                       // mm_interconnect_0:C3_s1_address -> C3:address
	wire  [31:0] mm_interconnect_0_c2_s1_readdata;                      // C2:readdata -> mm_interconnect_0:C2_s1_readdata
	wire   [1:0] mm_interconnect_0_c2_s1_address;                       // mm_interconnect_0:C2_s1_address -> C2:address
	wire  [31:0] mm_interconnect_0_c1_s1_readdata;                      // C1:readdata -> mm_interconnect_0:C1_s1_readdata
	wire   [1:0] mm_interconnect_0_c1_s1_address;                       // mm_interconnect_0:C1_s1_address -> C1:address
	wire         mm_interconnect_0_r4_s1_chipselect;                    // mm_interconnect_0:R4_s1_chipselect -> R4:chipselect
	wire  [31:0] mm_interconnect_0_r4_s1_readdata;                      // R4:readdata -> mm_interconnect_0:R4_s1_readdata
	wire   [1:0] mm_interconnect_0_r4_s1_address;                       // mm_interconnect_0:R4_s1_address -> R4:address
	wire         mm_interconnect_0_r4_s1_write;                         // mm_interconnect_0:R4_s1_write -> R4:write_n
	wire  [31:0] mm_interconnect_0_r4_s1_writedata;                     // mm_interconnect_0:R4_s1_writedata -> R4:writedata
	wire         mm_interconnect_0_r3_s1_chipselect;                    // mm_interconnect_0:R3_s1_chipselect -> R3:chipselect
	wire  [31:0] mm_interconnect_0_r3_s1_readdata;                      // R3:readdata -> mm_interconnect_0:R3_s1_readdata
	wire   [1:0] mm_interconnect_0_r3_s1_address;                       // mm_interconnect_0:R3_s1_address -> R3:address
	wire         mm_interconnect_0_r3_s1_write;                         // mm_interconnect_0:R3_s1_write -> R3:write_n
	wire  [31:0] mm_interconnect_0_r3_s1_writedata;                     // mm_interconnect_0:R3_s1_writedata -> R3:writedata
	wire         mm_interconnect_0_r2_s1_chipselect;                    // mm_interconnect_0:R2_s1_chipselect -> R2:chipselect
	wire  [31:0] mm_interconnect_0_r2_s1_readdata;                      // R2:readdata -> mm_interconnect_0:R2_s1_readdata
	wire   [1:0] mm_interconnect_0_r2_s1_address;                       // mm_interconnect_0:R2_s1_address -> R2:address
	wire         mm_interconnect_0_r2_s1_write;                         // mm_interconnect_0:R2_s1_write -> R2:write_n
	wire  [31:0] mm_interconnect_0_r2_s1_writedata;                     // mm_interconnect_0:R2_s1_writedata -> R2:writedata
	wire         mm_interconnect_0_r1_s1_chipselect;                    // mm_interconnect_0:R1_s1_chipselect -> R1:chipselect
	wire  [31:0] mm_interconnect_0_r1_s1_readdata;                      // R1:readdata -> mm_interconnect_0:R1_s1_readdata
	wire   [1:0] mm_interconnect_0_r1_s1_address;                       // mm_interconnect_0:R1_s1_address -> R1:address
	wire         mm_interconnect_0_r1_s1_write;                         // mm_interconnect_0:R1_s1_write -> R1:write_n
	wire  [31:0] mm_interconnect_0_r1_s1_writedata;                     // mm_interconnect_0:R1_s1_writedata -> R1:writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                   // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                     // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [15:0] mm_interconnect_0_ram_s1_address;                      // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                   // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                        // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                    // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                        // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         mm_interconnect_0_timer_0_s1_chipselect;               // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                 // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                  // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                    // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         irq_mapper_receiver0_irq;                              // DEBUG:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                              // timer_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_irq_irq;                                           // irq_mapper:sender_irq -> CPU:irq
	wire         rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [C1:reset_n, C2:reset_n, C3:reset_n, C4:reset_n, CPU:reset_n, DEBUG:rst_n, R1:reset_n, R2:reset_n, R3:reset_n, R4:reset_n, RAM:reset, irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset, rst_translator:in_reset, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                    // rst_controller:reset_req -> [CPU:reset_req, RAM:reset_req, rst_translator:reset_req_in]

	ledMatrix_C1 c1 (
		.clk      (clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_c1_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_c1_s1_readdata), //                    .readdata
		.in_port  (c1_export)                         // external_connection.export
	);

	ledMatrix_C1 c2 (
		.clk      (clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_c2_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_c2_s1_readdata), //                    .readdata
		.in_port  (c2_export)                         // external_connection.export
	);

	ledMatrix_C1 c3 (
		.clk      (clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_c3_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_c3_s1_readdata), //                    .readdata
		.in_port  (c3_export)                         // external_connection.export
	);

	ledMatrix_C1 c4 (
		.clk      (clk_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_c4_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_c4_s1_readdata), //                    .readdata
		.in_port  (c4_export)                         // external_connection.export
	);

	ledMatrix_CPU cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                  //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	ledMatrix_DEBUG debug (
		.clk            (clk_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_debug_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_debug_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_debug_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                               //               irq.irq
	);

	ledMatrix_R1 r1 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_r1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_r1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_r1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_r1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_r1_s1_readdata),   //                    .readdata
		.out_port   (r1_export)                           // external_connection.export
	);

	ledMatrix_R1 r2 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_r2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_r2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_r2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_r2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_r2_s1_readdata),   //                    .readdata
		.out_port   (r2_export)                           // external_connection.export
	);

	ledMatrix_R1 r3 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_r3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_r3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_r3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_r3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_r3_s1_readdata),   //                    .readdata
		.out_port   (r3_export)                           // external_connection.export
	);

	ledMatrix_R1 r4 (
		.clk        (clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),    //               reset.reset_n
		.address    (mm_interconnect_0_r4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_r4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_r4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_r4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_r4_s1_readdata),   //                    .readdata
		.out_port   (r4_export)                           // external_connection.export
	);

	ledMatrix_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	ledMatrix_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	ledMatrix_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                         (clk_clk),                                               //                       clk_0_clk.clk
		.CPU_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                        // CPU_reset_reset_bridge_in_reset.reset
		.CPU_data_master_address               (cpu_data_master_address),                               //                 CPU_data_master.address
		.CPU_data_master_waitrequest           (cpu_data_master_waitrequest),                           //                                .waitrequest
		.CPU_data_master_byteenable            (cpu_data_master_byteenable),                            //                                .byteenable
		.CPU_data_master_read                  (cpu_data_master_read),                                  //                                .read
		.CPU_data_master_readdata              (cpu_data_master_readdata),                              //                                .readdata
		.CPU_data_master_write                 (cpu_data_master_write),                                 //                                .write
		.CPU_data_master_writedata             (cpu_data_master_writedata),                             //                                .writedata
		.CPU_data_master_debugaccess           (cpu_data_master_debugaccess),                           //                                .debugaccess
		.CPU_instruction_master_address        (cpu_instruction_master_address),                        //          CPU_instruction_master.address
		.CPU_instruction_master_waitrequest    (cpu_instruction_master_waitrequest),                    //                                .waitrequest
		.CPU_instruction_master_read           (cpu_instruction_master_read),                           //                                .read
		.CPU_instruction_master_readdata       (cpu_instruction_master_readdata),                       //                                .readdata
		.C1_s1_address                         (mm_interconnect_0_c1_s1_address),                       //                           C1_s1.address
		.C1_s1_readdata                        (mm_interconnect_0_c1_s1_readdata),                      //                                .readdata
		.C2_s1_address                         (mm_interconnect_0_c2_s1_address),                       //                           C2_s1.address
		.C2_s1_readdata                        (mm_interconnect_0_c2_s1_readdata),                      //                                .readdata
		.C3_s1_address                         (mm_interconnect_0_c3_s1_address),                       //                           C3_s1.address
		.C3_s1_readdata                        (mm_interconnect_0_c3_s1_readdata),                      //                                .readdata
		.C4_s1_address                         (mm_interconnect_0_c4_s1_address),                       //                           C4_s1.address
		.C4_s1_readdata                        (mm_interconnect_0_c4_s1_readdata),                      //                                .readdata
		.CPU_debug_mem_slave_address           (mm_interconnect_0_cpu_debug_mem_slave_address),         //             CPU_debug_mem_slave.address
		.CPU_debug_mem_slave_write             (mm_interconnect_0_cpu_debug_mem_slave_write),           //                                .write
		.CPU_debug_mem_slave_read              (mm_interconnect_0_cpu_debug_mem_slave_read),            //                                .read
		.CPU_debug_mem_slave_readdata          (mm_interconnect_0_cpu_debug_mem_slave_readdata),        //                                .readdata
		.CPU_debug_mem_slave_writedata         (mm_interconnect_0_cpu_debug_mem_slave_writedata),       //                                .writedata
		.CPU_debug_mem_slave_byteenable        (mm_interconnect_0_cpu_debug_mem_slave_byteenable),      //                                .byteenable
		.CPU_debug_mem_slave_waitrequest       (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),     //                                .waitrequest
		.CPU_debug_mem_slave_debugaccess       (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),     //                                .debugaccess
		.DEBUG_avalon_jtag_slave_address       (mm_interconnect_0_debug_avalon_jtag_slave_address),     //         DEBUG_avalon_jtag_slave.address
		.DEBUG_avalon_jtag_slave_write         (mm_interconnect_0_debug_avalon_jtag_slave_write),       //                                .write
		.DEBUG_avalon_jtag_slave_read          (mm_interconnect_0_debug_avalon_jtag_slave_read),        //                                .read
		.DEBUG_avalon_jtag_slave_readdata      (mm_interconnect_0_debug_avalon_jtag_slave_readdata),    //                                .readdata
		.DEBUG_avalon_jtag_slave_writedata     (mm_interconnect_0_debug_avalon_jtag_slave_writedata),   //                                .writedata
		.DEBUG_avalon_jtag_slave_waitrequest   (mm_interconnect_0_debug_avalon_jtag_slave_waitrequest), //                                .waitrequest
		.DEBUG_avalon_jtag_slave_chipselect    (mm_interconnect_0_debug_avalon_jtag_slave_chipselect),  //                                .chipselect
		.R1_s1_address                         (mm_interconnect_0_r1_s1_address),                       //                           R1_s1.address
		.R1_s1_write                           (mm_interconnect_0_r1_s1_write),                         //                                .write
		.R1_s1_readdata                        (mm_interconnect_0_r1_s1_readdata),                      //                                .readdata
		.R1_s1_writedata                       (mm_interconnect_0_r1_s1_writedata),                     //                                .writedata
		.R1_s1_chipselect                      (mm_interconnect_0_r1_s1_chipselect),                    //                                .chipselect
		.R2_s1_address                         (mm_interconnect_0_r2_s1_address),                       //                           R2_s1.address
		.R2_s1_write                           (mm_interconnect_0_r2_s1_write),                         //                                .write
		.R2_s1_readdata                        (mm_interconnect_0_r2_s1_readdata),                      //                                .readdata
		.R2_s1_writedata                       (mm_interconnect_0_r2_s1_writedata),                     //                                .writedata
		.R2_s1_chipselect                      (mm_interconnect_0_r2_s1_chipselect),                    //                                .chipselect
		.R3_s1_address                         (mm_interconnect_0_r3_s1_address),                       //                           R3_s1.address
		.R3_s1_write                           (mm_interconnect_0_r3_s1_write),                         //                                .write
		.R3_s1_readdata                        (mm_interconnect_0_r3_s1_readdata),                      //                                .readdata
		.R3_s1_writedata                       (mm_interconnect_0_r3_s1_writedata),                     //                                .writedata
		.R3_s1_chipselect                      (mm_interconnect_0_r3_s1_chipselect),                    //                                .chipselect
		.R4_s1_address                         (mm_interconnect_0_r4_s1_address),                       //                           R4_s1.address
		.R4_s1_write                           (mm_interconnect_0_r4_s1_write),                         //                                .write
		.R4_s1_readdata                        (mm_interconnect_0_r4_s1_readdata),                      //                                .readdata
		.R4_s1_writedata                       (mm_interconnect_0_r4_s1_writedata),                     //                                .writedata
		.R4_s1_chipselect                      (mm_interconnect_0_r4_s1_chipselect),                    //                                .chipselect
		.RAM_s1_address                        (mm_interconnect_0_ram_s1_address),                      //                          RAM_s1.address
		.RAM_s1_write                          (mm_interconnect_0_ram_s1_write),                        //                                .write
		.RAM_s1_readdata                       (mm_interconnect_0_ram_s1_readdata),                     //                                .readdata
		.RAM_s1_writedata                      (mm_interconnect_0_ram_s1_writedata),                    //                                .writedata
		.RAM_s1_byteenable                     (mm_interconnect_0_ram_s1_byteenable),                   //                                .byteenable
		.RAM_s1_chipselect                     (mm_interconnect_0_ram_s1_chipselect),                   //                                .chipselect
		.RAM_s1_clken                          (mm_interconnect_0_ram_s1_clken),                        //                                .clken
		.timer_0_s1_address                    (mm_interconnect_0_timer_0_s1_address),                  //                      timer_0_s1.address
		.timer_0_s1_write                      (mm_interconnect_0_timer_0_s1_write),                    //                                .write
		.timer_0_s1_readdata                   (mm_interconnect_0_timer_0_s1_readdata),                 //                                .readdata
		.timer_0_s1_writedata                  (mm_interconnect_0_timer_0_s1_writedata),                //                                .writedata
		.timer_0_s1_chipselect                 (mm_interconnect_0_timer_0_s1_chipselect)                //                                .chipselect
	);

	ledMatrix_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
