
module interrupt (
	clk_clk,
	reset_reset_n,
	led_export,
	button_export);	

	input		clk_clk;
	input		reset_reset_n;
	output		led_export;
	input		button_export;
endmodule
