// sdram.v

// Generated using ACDS version 22.1 915

`timescale 1 ps / 1 ps
module sdram (
		output wire        aux_full_rate_clk,  // aux_full_rate_clk.clk
		output wire        aux_half_rate_clk,  // aux_half_rate_clk.clk
		output wire        local_ready,        //               avl.waitrequest_n
		input  wire        local_write_req,    //                  .write
		input  wire        local_read_req,     //                  .read
		input  wire [23:0] local_address,      //                  .address
		input  wire [1:0]  local_be,           //                  .byteenable
		input  wire [15:0] local_wdata,        //                  .writedata
		input  wire [2:0]  local_size,         //                  .burstcount
		input  wire        local_burstbegin,   //                  .beginbursttransfer
		output wire [15:0] local_rdata,        //                  .readdata
		output wire        local_rdata_valid,  //                  .readdatavalid
		input  wire        global_reset_n,     //      global_reset.reset_n
		output wire [12:0] mem_addr,           //               mem.mem_a
		output wire [1:0]  mem_ba,             //                  .mem_ba
		output wire        mem_cas_n,          //                  .mem_cas_n
		output wire        mem_cke,            //                  .mem_cke
		inout  wire        mem_clk,            //                  .mem_ck
		inout  wire        mem_clk_n,          //                  .mem_ck_n
		output wire        mem_cs_n,           //                  .mem_cs_n
		output wire        mem_dm,             //                  .mem_dm
		inout  wire [7:0]  mem_dq,             //                  .mem_dq
		inout  wire        mem_dqs,            //                  .mem_dqs
		inout  wire        mem_dqs_n,          //                  .mem_dqs_n
		output wire        mem_odt,            //                  .mem_odt
		output wire        mem_ras_n,          //                  .mem_ras_n
		output wire        mem_we_n,           //                  .mem_we_n
		output wire        phy_clk,            //           phy_clk.clk
		output wire        reset_phy_clk_n,    //         phy_reset.reset_n
		input  wire        pll_ref_clk,        //       pll_ref_clk.clk
		output wire        reset_request_n,    //     reset_request.reset_n
		output wire        status_cal_fail,    //            status.local_cal_fail
		output wire        status_cal_success, //                  .local_cal_success
		output wire        status_init_done    //                  .local_init_done
	);

	sdram_alt_mem_if_civ_ddr2_emif_0 alt_mem_if_civ_ddr2_emif_0 (
		.phy_clk            (phy_clk),            //           phy_clk.clk
		.reset_phy_clk_n    (reset_phy_clk_n),    //         phy_reset.reset_n
		.status_cal_fail    (status_cal_fail),    //            status.local_cal_fail
		.status_cal_success (status_cal_success), //                  .local_cal_success
		.status_init_done   (status_init_done),   //                  .local_init_done
		.global_reset_n     (global_reset_n),     //      global_reset.reset_n
		.reset_request_n    (reset_request_n),    //     reset_request.reset_n
		.local_ready        (local_ready),        //               avl.waitrequest_n
		.local_write_req    (local_write_req),    //                  .write
		.local_read_req     (local_read_req),     //                  .read
		.local_address      (local_address),      //                  .address
		.local_be           (local_be),           //                  .byteenable
		.local_wdata        (local_wdata),        //                  .writedata
		.local_size         (local_size),         //                  .burstcount
		.local_burstbegin   (local_burstbegin),   //                  .beginbursttransfer
		.local_rdata        (local_rdata),        //                  .readdata
		.local_rdata_valid  (local_rdata_valid),  //                  .readdatavalid
		.mem_addr           (mem_addr),           //               mem.mem_a
		.mem_ba             (mem_ba),             //                  .mem_ba
		.mem_cas_n          (mem_cas_n),          //                  .mem_cas_n
		.mem_cke            (mem_cke),            //                  .mem_cke
		.mem_clk            (mem_clk),            //                  .mem_ck
		.mem_clk_n          (mem_clk_n),          //                  .mem_ck_n
		.mem_cs_n           (mem_cs_n),           //                  .mem_cs_n
		.mem_dm             (mem_dm),             //                  .mem_dm
		.mem_dq             (mem_dq),             //                  .mem_dq
		.mem_dqs            (mem_dqs),            //                  .mem_dqs
		.mem_dqs_n          (mem_dqs_n),          //                  .mem_dqs_n
		.mem_odt            (mem_odt),            //                  .mem_odt
		.mem_ras_n          (mem_ras_n),          //                  .mem_ras_n
		.mem_we_n           (mem_we_n),           //                  .mem_we_n
		.aux_full_rate_clk  (aux_full_rate_clk),  // aux_full_rate_clk.clk
		.aux_half_rate_clk  (aux_half_rate_clk),  // aux_half_rate_clk.clk
		.pll_ref_clk        (pll_ref_clk)         //       pll_ref_clk.clk
	);

endmodule
